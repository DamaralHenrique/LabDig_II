-- Calibrador + registradores